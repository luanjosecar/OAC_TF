-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_MUX 

-- ============================================================
-- File Name: mux324.vhd
-- Megafunction Name(s):
-- 			LPM_MUX
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY mux324 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data16x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data17x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data18x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data19x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data20x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data21x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data22x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data23x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data24x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data25x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data26x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data27x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data28x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data29x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data30x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data31x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END mux324;


ARCHITECTURE SYN OF mux324 IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_2D (31 DOWNTO 0, 31 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire18	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire19	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire20	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire21	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire22	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire23	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire24	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire25	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire26	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire27	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire28	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire29	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire30	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire31	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire32	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire33	: STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
	sub_wire33    <= data0x(31 DOWNTO 0);
	sub_wire32    <= data1x(31 DOWNTO 0);
	sub_wire31    <= data2x(31 DOWNTO 0);
	sub_wire30    <= data3x(31 DOWNTO 0);
	sub_wire29    <= data4x(31 DOWNTO 0);
	sub_wire28    <= data5x(31 DOWNTO 0);
	sub_wire27    <= data6x(31 DOWNTO 0);
	sub_wire26    <= data7x(31 DOWNTO 0);
	sub_wire25    <= data8x(31 DOWNTO 0);
	sub_wire24    <= data9x(31 DOWNTO 0);
	sub_wire23    <= data10x(31 DOWNTO 0);
	sub_wire22    <= data11x(31 DOWNTO 0);
	sub_wire21    <= data12x(31 DOWNTO 0);
	sub_wire20    <= data13x(31 DOWNTO 0);
	sub_wire19    <= data14x(31 DOWNTO 0);
	sub_wire18    <= data15x(31 DOWNTO 0);
	sub_wire17    <= data16x(31 DOWNTO 0);
	sub_wire16    <= data17x(31 DOWNTO 0);
	sub_wire15    <= data18x(31 DOWNTO 0);
	sub_wire14    <= data19x(31 DOWNTO 0);
	sub_wire13    <= data20x(31 DOWNTO 0);
	sub_wire12    <= data21x(31 DOWNTO 0);
	sub_wire11    <= data22x(31 DOWNTO 0);
	sub_wire10    <= data23x(31 DOWNTO 0);
	sub_wire9    <= data24x(31 DOWNTO 0);
	sub_wire8    <= data25x(31 DOWNTO 0);
	sub_wire7    <= data26x(31 DOWNTO 0);
	sub_wire6    <= data27x(31 DOWNTO 0);
	sub_wire5    <= data28x(31 DOWNTO 0);
	sub_wire4    <= data29x(31 DOWNTO 0);
	sub_wire3    <= data30x(31 DOWNTO 0);
	result    <= sub_wire0(31 DOWNTO 0);
	sub_wire1    <= data31x(31 DOWNTO 0);
	sub_wire2(31, 0)    <= sub_wire1(0);
	sub_wire2(31, 1)    <= sub_wire1(1);
	sub_wire2(31, 2)    <= sub_wire1(2);
	sub_wire2(31, 3)    <= sub_wire1(3);
	sub_wire2(31, 4)    <= sub_wire1(4);
	sub_wire2(31, 5)    <= sub_wire1(5);
	sub_wire2(31, 6)    <= sub_wire1(6);
	sub_wire2(31, 7)    <= sub_wire1(7);
	sub_wire2(31, 8)    <= sub_wire1(8);
	sub_wire2(31, 9)    <= sub_wire1(9);
	sub_wire2(31, 10)    <= sub_wire1(10);
	sub_wire2(31, 11)    <= sub_wire1(11);
	sub_wire2(31, 12)    <= sub_wire1(12);
	sub_wire2(31, 13)    <= sub_wire1(13);
	sub_wire2(31, 14)    <= sub_wire1(14);
	sub_wire2(31, 15)    <= sub_wire1(15);
	sub_wire2(31, 16)    <= sub_wire1(16);
	sub_wire2(31, 17)    <= sub_wire1(17);
	sub_wire2(31, 18)    <= sub_wire1(18);
	sub_wire2(31, 19)    <= sub_wire1(19);
	sub_wire2(31, 20)    <= sub_wire1(20);
	sub_wire2(31, 21)    <= sub_wire1(21);
	sub_wire2(31, 22)    <= sub_wire1(22);
	sub_wire2(31, 23)    <= sub_wire1(23);
	sub_wire2(31, 24)    <= sub_wire1(24);
	sub_wire2(31, 25)    <= sub_wire1(25);
	sub_wire2(31, 26)    <= sub_wire1(26);
	sub_wire2(31, 27)    <= sub_wire1(27);
	sub_wire2(31, 28)    <= sub_wire1(28);
	sub_wire2(31, 29)    <= sub_wire1(29);
	sub_wire2(31, 30)    <= sub_wire1(30);
	sub_wire2(31, 31)    <= sub_wire1(31);
	sub_wire2(30, 0)    <= sub_wire3(0);
	sub_wire2(30, 1)    <= sub_wire3(1);
	sub_wire2(30, 2)    <= sub_wire3(2);
	sub_wire2(30, 3)    <= sub_wire3(3);
	sub_wire2(30, 4)    <= sub_wire3(4);
	sub_wire2(30, 5)    <= sub_wire3(5);
	sub_wire2(30, 6)    <= sub_wire3(6);
	sub_wire2(30, 7)    <= sub_wire3(7);
	sub_wire2(30, 8)    <= sub_wire3(8);
	sub_wire2(30, 9)    <= sub_wire3(9);
	sub_wire2(30, 10)    <= sub_wire3(10);
	sub_wire2(30, 11)    <= sub_wire3(11);
	sub_wire2(30, 12)    <= sub_wire3(12);
	sub_wire2(30, 13)    <= sub_wire3(13);
	sub_wire2(30, 14)    <= sub_wire3(14);
	sub_wire2(30, 15)    <= sub_wire3(15);
	sub_wire2(30, 16)    <= sub_wire3(16);
	sub_wire2(30, 17)    <= sub_wire3(17);
	sub_wire2(30, 18)    <= sub_wire3(18);
	sub_wire2(30, 19)    <= sub_wire3(19);
	sub_wire2(30, 20)    <= sub_wire3(20);
	sub_wire2(30, 21)    <= sub_wire3(21);
	sub_wire2(30, 22)    <= sub_wire3(22);
	sub_wire2(30, 23)    <= sub_wire3(23);
	sub_wire2(30, 24)    <= sub_wire3(24);
	sub_wire2(30, 25)    <= sub_wire3(25);
	sub_wire2(30, 26)    <= sub_wire3(26);
	sub_wire2(30, 27)    <= sub_wire3(27);
	sub_wire2(30, 28)    <= sub_wire3(28);
	sub_wire2(30, 29)    <= sub_wire3(29);
	sub_wire2(30, 30)    <= sub_wire3(30);
	sub_wire2(30, 31)    <= sub_wire3(31);
	sub_wire2(29, 0)    <= sub_wire4(0);
	sub_wire2(29, 1)    <= sub_wire4(1);
	sub_wire2(29, 2)    <= sub_wire4(2);
	sub_wire2(29, 3)    <= sub_wire4(3);
	sub_wire2(29, 4)    <= sub_wire4(4);
	sub_wire2(29, 5)    <= sub_wire4(5);
	sub_wire2(29, 6)    <= sub_wire4(6);
	sub_wire2(29, 7)    <= sub_wire4(7);
	sub_wire2(29, 8)    <= sub_wire4(8);
	sub_wire2(29, 9)    <= sub_wire4(9);
	sub_wire2(29, 10)    <= sub_wire4(10);
	sub_wire2(29, 11)    <= sub_wire4(11);
	sub_wire2(29, 12)    <= sub_wire4(12);
	sub_wire2(29, 13)    <= sub_wire4(13);
	sub_wire2(29, 14)    <= sub_wire4(14);
	sub_wire2(29, 15)    <= sub_wire4(15);
	sub_wire2(29, 16)    <= sub_wire4(16);
	sub_wire2(29, 17)    <= sub_wire4(17);
	sub_wire2(29, 18)    <= sub_wire4(18);
	sub_wire2(29, 19)    <= sub_wire4(19);
	sub_wire2(29, 20)    <= sub_wire4(20);
	sub_wire2(29, 21)    <= sub_wire4(21);
	sub_wire2(29, 22)    <= sub_wire4(22);
	sub_wire2(29, 23)    <= sub_wire4(23);
	sub_wire2(29, 24)    <= sub_wire4(24);
	sub_wire2(29, 25)    <= sub_wire4(25);
	sub_wire2(29, 26)    <= sub_wire4(26);
	sub_wire2(29, 27)    <= sub_wire4(27);
	sub_wire2(29, 28)    <= sub_wire4(28);
	sub_wire2(29, 29)    <= sub_wire4(29);
	sub_wire2(29, 30)    <= sub_wire4(30);
	sub_wire2(29, 31)    <= sub_wire4(31);
	sub_wire2(28, 0)    <= sub_wire5(0);
	sub_wire2(28, 1)    <= sub_wire5(1);
	sub_wire2(28, 2)    <= sub_wire5(2);
	sub_wire2(28, 3)    <= sub_wire5(3);
	sub_wire2(28, 4)    <= sub_wire5(4);
	sub_wire2(28, 5)    <= sub_wire5(5);
	sub_wire2(28, 6)    <= sub_wire5(6);
	sub_wire2(28, 7)    <= sub_wire5(7);
	sub_wire2(28, 8)    <= sub_wire5(8);
	sub_wire2(28, 9)    <= sub_wire5(9);
	sub_wire2(28, 10)    <= sub_wire5(10);
	sub_wire2(28, 11)    <= sub_wire5(11);
	sub_wire2(28, 12)    <= sub_wire5(12);
	sub_wire2(28, 13)    <= sub_wire5(13);
	sub_wire2(28, 14)    <= sub_wire5(14);
	sub_wire2(28, 15)    <= sub_wire5(15);
	sub_wire2(28, 16)    <= sub_wire5(16);
	sub_wire2(28, 17)    <= sub_wire5(17);
	sub_wire2(28, 18)    <= sub_wire5(18);
	sub_wire2(28, 19)    <= sub_wire5(19);
	sub_wire2(28, 20)    <= sub_wire5(20);
	sub_wire2(28, 21)    <= sub_wire5(21);
	sub_wire2(28, 22)    <= sub_wire5(22);
	sub_wire2(28, 23)    <= sub_wire5(23);
	sub_wire2(28, 24)    <= sub_wire5(24);
	sub_wire2(28, 25)    <= sub_wire5(25);
	sub_wire2(28, 26)    <= sub_wire5(26);
	sub_wire2(28, 27)    <= sub_wire5(27);
	sub_wire2(28, 28)    <= sub_wire5(28);
	sub_wire2(28, 29)    <= sub_wire5(29);
	sub_wire2(28, 30)    <= sub_wire5(30);
	sub_wire2(28, 31)    <= sub_wire5(31);
	sub_wire2(27, 0)    <= sub_wire6(0);
	sub_wire2(27, 1)    <= sub_wire6(1);
	sub_wire2(27, 2)    <= sub_wire6(2);
	sub_wire2(27, 3)    <= sub_wire6(3);
	sub_wire2(27, 4)    <= sub_wire6(4);
	sub_wire2(27, 5)    <= sub_wire6(5);
	sub_wire2(27, 6)    <= sub_wire6(6);
	sub_wire2(27, 7)    <= sub_wire6(7);
	sub_wire2(27, 8)    <= sub_wire6(8);
	sub_wire2(27, 9)    <= sub_wire6(9);
	sub_wire2(27, 10)    <= sub_wire6(10);
	sub_wire2(27, 11)    <= sub_wire6(11);
	sub_wire2(27, 12)    <= sub_wire6(12);
	sub_wire2(27, 13)    <= sub_wire6(13);
	sub_wire2(27, 14)    <= sub_wire6(14);
	sub_wire2(27, 15)    <= sub_wire6(15);
	sub_wire2(27, 16)    <= sub_wire6(16);
	sub_wire2(27, 17)    <= sub_wire6(17);
	sub_wire2(27, 18)    <= sub_wire6(18);
	sub_wire2(27, 19)    <= sub_wire6(19);
	sub_wire2(27, 20)    <= sub_wire6(20);
	sub_wire2(27, 21)    <= sub_wire6(21);
	sub_wire2(27, 22)    <= sub_wire6(22);
	sub_wire2(27, 23)    <= sub_wire6(23);
	sub_wire2(27, 24)    <= sub_wire6(24);
	sub_wire2(27, 25)    <= sub_wire6(25);
	sub_wire2(27, 26)    <= sub_wire6(26);
	sub_wire2(27, 27)    <= sub_wire6(27);
	sub_wire2(27, 28)    <= sub_wire6(28);
	sub_wire2(27, 29)    <= sub_wire6(29);
	sub_wire2(27, 30)    <= sub_wire6(30);
	sub_wire2(27, 31)    <= sub_wire6(31);
	sub_wire2(26, 0)    <= sub_wire7(0);
	sub_wire2(26, 1)    <= sub_wire7(1);
	sub_wire2(26, 2)    <= sub_wire7(2);
	sub_wire2(26, 3)    <= sub_wire7(3);
	sub_wire2(26, 4)    <= sub_wire7(4);
	sub_wire2(26, 5)    <= sub_wire7(5);
	sub_wire2(26, 6)    <= sub_wire7(6);
	sub_wire2(26, 7)    <= sub_wire7(7);
	sub_wire2(26, 8)    <= sub_wire7(8);
	sub_wire2(26, 9)    <= sub_wire7(9);
	sub_wire2(26, 10)    <= sub_wire7(10);
	sub_wire2(26, 11)    <= sub_wire7(11);
	sub_wire2(26, 12)    <= sub_wire7(12);
	sub_wire2(26, 13)    <= sub_wire7(13);
	sub_wire2(26, 14)    <= sub_wire7(14);
	sub_wire2(26, 15)    <= sub_wire7(15);
	sub_wire2(26, 16)    <= sub_wire7(16);
	sub_wire2(26, 17)    <= sub_wire7(17);
	sub_wire2(26, 18)    <= sub_wire7(18);
	sub_wire2(26, 19)    <= sub_wire7(19);
	sub_wire2(26, 20)    <= sub_wire7(20);
	sub_wire2(26, 21)    <= sub_wire7(21);
	sub_wire2(26, 22)    <= sub_wire7(22);
	sub_wire2(26, 23)    <= sub_wire7(23);
	sub_wire2(26, 24)    <= sub_wire7(24);
	sub_wire2(26, 25)    <= sub_wire7(25);
	sub_wire2(26, 26)    <= sub_wire7(26);
	sub_wire2(26, 27)    <= sub_wire7(27);
	sub_wire2(26, 28)    <= sub_wire7(28);
	sub_wire2(26, 29)    <= sub_wire7(29);
	sub_wire2(26, 30)    <= sub_wire7(30);
	sub_wire2(26, 31)    <= sub_wire7(31);
	sub_wire2(25, 0)    <= sub_wire8(0);
	sub_wire2(25, 1)    <= sub_wire8(1);
	sub_wire2(25, 2)    <= sub_wire8(2);
	sub_wire2(25, 3)    <= sub_wire8(3);
	sub_wire2(25, 4)    <= sub_wire8(4);
	sub_wire2(25, 5)    <= sub_wire8(5);
	sub_wire2(25, 6)    <= sub_wire8(6);
	sub_wire2(25, 7)    <= sub_wire8(7);
	sub_wire2(25, 8)    <= sub_wire8(8);
	sub_wire2(25, 9)    <= sub_wire8(9);
	sub_wire2(25, 10)    <= sub_wire8(10);
	sub_wire2(25, 11)    <= sub_wire8(11);
	sub_wire2(25, 12)    <= sub_wire8(12);
	sub_wire2(25, 13)    <= sub_wire8(13);
	sub_wire2(25, 14)    <= sub_wire8(14);
	sub_wire2(25, 15)    <= sub_wire8(15);
	sub_wire2(25, 16)    <= sub_wire8(16);
	sub_wire2(25, 17)    <= sub_wire8(17);
	sub_wire2(25, 18)    <= sub_wire8(18);
	sub_wire2(25, 19)    <= sub_wire8(19);
	sub_wire2(25, 20)    <= sub_wire8(20);
	sub_wire2(25, 21)    <= sub_wire8(21);
	sub_wire2(25, 22)    <= sub_wire8(22);
	sub_wire2(25, 23)    <= sub_wire8(23);
	sub_wire2(25, 24)    <= sub_wire8(24);
	sub_wire2(25, 25)    <= sub_wire8(25);
	sub_wire2(25, 26)    <= sub_wire8(26);
	sub_wire2(25, 27)    <= sub_wire8(27);
	sub_wire2(25, 28)    <= sub_wire8(28);
	sub_wire2(25, 29)    <= sub_wire8(29);
	sub_wire2(25, 30)    <= sub_wire8(30);
	sub_wire2(25, 31)    <= sub_wire8(31);
	sub_wire2(24, 0)    <= sub_wire9(0);
	sub_wire2(24, 1)    <= sub_wire9(1);
	sub_wire2(24, 2)    <= sub_wire9(2);
	sub_wire2(24, 3)    <= sub_wire9(3);
	sub_wire2(24, 4)    <= sub_wire9(4);
	sub_wire2(24, 5)    <= sub_wire9(5);
	sub_wire2(24, 6)    <= sub_wire9(6);
	sub_wire2(24, 7)    <= sub_wire9(7);
	sub_wire2(24, 8)    <= sub_wire9(8);
	sub_wire2(24, 9)    <= sub_wire9(9);
	sub_wire2(24, 10)    <= sub_wire9(10);
	sub_wire2(24, 11)    <= sub_wire9(11);
	sub_wire2(24, 12)    <= sub_wire9(12);
	sub_wire2(24, 13)    <= sub_wire9(13);
	sub_wire2(24, 14)    <= sub_wire9(14);
	sub_wire2(24, 15)    <= sub_wire9(15);
	sub_wire2(24, 16)    <= sub_wire9(16);
	sub_wire2(24, 17)    <= sub_wire9(17);
	sub_wire2(24, 18)    <= sub_wire9(18);
	sub_wire2(24, 19)    <= sub_wire9(19);
	sub_wire2(24, 20)    <= sub_wire9(20);
	sub_wire2(24, 21)    <= sub_wire9(21);
	sub_wire2(24, 22)    <= sub_wire9(22);
	sub_wire2(24, 23)    <= sub_wire9(23);
	sub_wire2(24, 24)    <= sub_wire9(24);
	sub_wire2(24, 25)    <= sub_wire9(25);
	sub_wire2(24, 26)    <= sub_wire9(26);
	sub_wire2(24, 27)    <= sub_wire9(27);
	sub_wire2(24, 28)    <= sub_wire9(28);
	sub_wire2(24, 29)    <= sub_wire9(29);
	sub_wire2(24, 30)    <= sub_wire9(30);
	sub_wire2(24, 31)    <= sub_wire9(31);
	sub_wire2(23, 0)    <= sub_wire10(0);
	sub_wire2(23, 1)    <= sub_wire10(1);
	sub_wire2(23, 2)    <= sub_wire10(2);
	sub_wire2(23, 3)    <= sub_wire10(3);
	sub_wire2(23, 4)    <= sub_wire10(4);
	sub_wire2(23, 5)    <= sub_wire10(5);
	sub_wire2(23, 6)    <= sub_wire10(6);
	sub_wire2(23, 7)    <= sub_wire10(7);
	sub_wire2(23, 8)    <= sub_wire10(8);
	sub_wire2(23, 9)    <= sub_wire10(9);
	sub_wire2(23, 10)    <= sub_wire10(10);
	sub_wire2(23, 11)    <= sub_wire10(11);
	sub_wire2(23, 12)    <= sub_wire10(12);
	sub_wire2(23, 13)    <= sub_wire10(13);
	sub_wire2(23, 14)    <= sub_wire10(14);
	sub_wire2(23, 15)    <= sub_wire10(15);
	sub_wire2(23, 16)    <= sub_wire10(16);
	sub_wire2(23, 17)    <= sub_wire10(17);
	sub_wire2(23, 18)    <= sub_wire10(18);
	sub_wire2(23, 19)    <= sub_wire10(19);
	sub_wire2(23, 20)    <= sub_wire10(20);
	sub_wire2(23, 21)    <= sub_wire10(21);
	sub_wire2(23, 22)    <= sub_wire10(22);
	sub_wire2(23, 23)    <= sub_wire10(23);
	sub_wire2(23, 24)    <= sub_wire10(24);
	sub_wire2(23, 25)    <= sub_wire10(25);
	sub_wire2(23, 26)    <= sub_wire10(26);
	sub_wire2(23, 27)    <= sub_wire10(27);
	sub_wire2(23, 28)    <= sub_wire10(28);
	sub_wire2(23, 29)    <= sub_wire10(29);
	sub_wire2(23, 30)    <= sub_wire10(30);
	sub_wire2(23, 31)    <= sub_wire10(31);
	sub_wire2(22, 0)    <= sub_wire11(0);
	sub_wire2(22, 1)    <= sub_wire11(1);
	sub_wire2(22, 2)    <= sub_wire11(2);
	sub_wire2(22, 3)    <= sub_wire11(3);
	sub_wire2(22, 4)    <= sub_wire11(4);
	sub_wire2(22, 5)    <= sub_wire11(5);
	sub_wire2(22, 6)    <= sub_wire11(6);
	sub_wire2(22, 7)    <= sub_wire11(7);
	sub_wire2(22, 8)    <= sub_wire11(8);
	sub_wire2(22, 9)    <= sub_wire11(9);
	sub_wire2(22, 10)    <= sub_wire11(10);
	sub_wire2(22, 11)    <= sub_wire11(11);
	sub_wire2(22, 12)    <= sub_wire11(12);
	sub_wire2(22, 13)    <= sub_wire11(13);
	sub_wire2(22, 14)    <= sub_wire11(14);
	sub_wire2(22, 15)    <= sub_wire11(15);
	sub_wire2(22, 16)    <= sub_wire11(16);
	sub_wire2(22, 17)    <= sub_wire11(17);
	sub_wire2(22, 18)    <= sub_wire11(18);
	sub_wire2(22, 19)    <= sub_wire11(19);
	sub_wire2(22, 20)    <= sub_wire11(20);
	sub_wire2(22, 21)    <= sub_wire11(21);
	sub_wire2(22, 22)    <= sub_wire11(22);
	sub_wire2(22, 23)    <= sub_wire11(23);
	sub_wire2(22, 24)    <= sub_wire11(24);
	sub_wire2(22, 25)    <= sub_wire11(25);
	sub_wire2(22, 26)    <= sub_wire11(26);
	sub_wire2(22, 27)    <= sub_wire11(27);
	sub_wire2(22, 28)    <= sub_wire11(28);
	sub_wire2(22, 29)    <= sub_wire11(29);
	sub_wire2(22, 30)    <= sub_wire11(30);
	sub_wire2(22, 31)    <= sub_wire11(31);
	sub_wire2(21, 0)    <= sub_wire12(0);
	sub_wire2(21, 1)    <= sub_wire12(1);
	sub_wire2(21, 2)    <= sub_wire12(2);
	sub_wire2(21, 3)    <= sub_wire12(3);
	sub_wire2(21, 4)    <= sub_wire12(4);
	sub_wire2(21, 5)    <= sub_wire12(5);
	sub_wire2(21, 6)    <= sub_wire12(6);
	sub_wire2(21, 7)    <= sub_wire12(7);
	sub_wire2(21, 8)    <= sub_wire12(8);
	sub_wire2(21, 9)    <= sub_wire12(9);
	sub_wire2(21, 10)    <= sub_wire12(10);
	sub_wire2(21, 11)    <= sub_wire12(11);
	sub_wire2(21, 12)    <= sub_wire12(12);
	sub_wire2(21, 13)    <= sub_wire12(13);
	sub_wire2(21, 14)    <= sub_wire12(14);
	sub_wire2(21, 15)    <= sub_wire12(15);
	sub_wire2(21, 16)    <= sub_wire12(16);
	sub_wire2(21, 17)    <= sub_wire12(17);
	sub_wire2(21, 18)    <= sub_wire12(18);
	sub_wire2(21, 19)    <= sub_wire12(19);
	sub_wire2(21, 20)    <= sub_wire12(20);
	sub_wire2(21, 21)    <= sub_wire12(21);
	sub_wire2(21, 22)    <= sub_wire12(22);
	sub_wire2(21, 23)    <= sub_wire12(23);
	sub_wire2(21, 24)    <= sub_wire12(24);
	sub_wire2(21, 25)    <= sub_wire12(25);
	sub_wire2(21, 26)    <= sub_wire12(26);
	sub_wire2(21, 27)    <= sub_wire12(27);
	sub_wire2(21, 28)    <= sub_wire12(28);
	sub_wire2(21, 29)    <= sub_wire12(29);
	sub_wire2(21, 30)    <= sub_wire12(30);
	sub_wire2(21, 31)    <= sub_wire12(31);
	sub_wire2(20, 0)    <= sub_wire13(0);
	sub_wire2(20, 1)    <= sub_wire13(1);
	sub_wire2(20, 2)    <= sub_wire13(2);
	sub_wire2(20, 3)    <= sub_wire13(3);
	sub_wire2(20, 4)    <= sub_wire13(4);
	sub_wire2(20, 5)    <= sub_wire13(5);
	sub_wire2(20, 6)    <= sub_wire13(6);
	sub_wire2(20, 7)    <= sub_wire13(7);
	sub_wire2(20, 8)    <= sub_wire13(8);
	sub_wire2(20, 9)    <= sub_wire13(9);
	sub_wire2(20, 10)    <= sub_wire13(10);
	sub_wire2(20, 11)    <= sub_wire13(11);
	sub_wire2(20, 12)    <= sub_wire13(12);
	sub_wire2(20, 13)    <= sub_wire13(13);
	sub_wire2(20, 14)    <= sub_wire13(14);
	sub_wire2(20, 15)    <= sub_wire13(15);
	sub_wire2(20, 16)    <= sub_wire13(16);
	sub_wire2(20, 17)    <= sub_wire13(17);
	sub_wire2(20, 18)    <= sub_wire13(18);
	sub_wire2(20, 19)    <= sub_wire13(19);
	sub_wire2(20, 20)    <= sub_wire13(20);
	sub_wire2(20, 21)    <= sub_wire13(21);
	sub_wire2(20, 22)    <= sub_wire13(22);
	sub_wire2(20, 23)    <= sub_wire13(23);
	sub_wire2(20, 24)    <= sub_wire13(24);
	sub_wire2(20, 25)    <= sub_wire13(25);
	sub_wire2(20, 26)    <= sub_wire13(26);
	sub_wire2(20, 27)    <= sub_wire13(27);
	sub_wire2(20, 28)    <= sub_wire13(28);
	sub_wire2(20, 29)    <= sub_wire13(29);
	sub_wire2(20, 30)    <= sub_wire13(30);
	sub_wire2(20, 31)    <= sub_wire13(31);
	sub_wire2(19, 0)    <= sub_wire14(0);
	sub_wire2(19, 1)    <= sub_wire14(1);
	sub_wire2(19, 2)    <= sub_wire14(2);
	sub_wire2(19, 3)    <= sub_wire14(3);
	sub_wire2(19, 4)    <= sub_wire14(4);
	sub_wire2(19, 5)    <= sub_wire14(5);
	sub_wire2(19, 6)    <= sub_wire14(6);
	sub_wire2(19, 7)    <= sub_wire14(7);
	sub_wire2(19, 8)    <= sub_wire14(8);
	sub_wire2(19, 9)    <= sub_wire14(9);
	sub_wire2(19, 10)    <= sub_wire14(10);
	sub_wire2(19, 11)    <= sub_wire14(11);
	sub_wire2(19, 12)    <= sub_wire14(12);
	sub_wire2(19, 13)    <= sub_wire14(13);
	sub_wire2(19, 14)    <= sub_wire14(14);
	sub_wire2(19, 15)    <= sub_wire14(15);
	sub_wire2(19, 16)    <= sub_wire14(16);
	sub_wire2(19, 17)    <= sub_wire14(17);
	sub_wire2(19, 18)    <= sub_wire14(18);
	sub_wire2(19, 19)    <= sub_wire14(19);
	sub_wire2(19, 20)    <= sub_wire14(20);
	sub_wire2(19, 21)    <= sub_wire14(21);
	sub_wire2(19, 22)    <= sub_wire14(22);
	sub_wire2(19, 23)    <= sub_wire14(23);
	sub_wire2(19, 24)    <= sub_wire14(24);
	sub_wire2(19, 25)    <= sub_wire14(25);
	sub_wire2(19, 26)    <= sub_wire14(26);
	sub_wire2(19, 27)    <= sub_wire14(27);
	sub_wire2(19, 28)    <= sub_wire14(28);
	sub_wire2(19, 29)    <= sub_wire14(29);
	sub_wire2(19, 30)    <= sub_wire14(30);
	sub_wire2(19, 31)    <= sub_wire14(31);
	sub_wire2(18, 0)    <= sub_wire15(0);
	sub_wire2(18, 1)    <= sub_wire15(1);
	sub_wire2(18, 2)    <= sub_wire15(2);
	sub_wire2(18, 3)    <= sub_wire15(3);
	sub_wire2(18, 4)    <= sub_wire15(4);
	sub_wire2(18, 5)    <= sub_wire15(5);
	sub_wire2(18, 6)    <= sub_wire15(6);
	sub_wire2(18, 7)    <= sub_wire15(7);
	sub_wire2(18, 8)    <= sub_wire15(8);
	sub_wire2(18, 9)    <= sub_wire15(9);
	sub_wire2(18, 10)    <= sub_wire15(10);
	sub_wire2(18, 11)    <= sub_wire15(11);
	sub_wire2(18, 12)    <= sub_wire15(12);
	sub_wire2(18, 13)    <= sub_wire15(13);
	sub_wire2(18, 14)    <= sub_wire15(14);
	sub_wire2(18, 15)    <= sub_wire15(15);
	sub_wire2(18, 16)    <= sub_wire15(16);
	sub_wire2(18, 17)    <= sub_wire15(17);
	sub_wire2(18, 18)    <= sub_wire15(18);
	sub_wire2(18, 19)    <= sub_wire15(19);
	sub_wire2(18, 20)    <= sub_wire15(20);
	sub_wire2(18, 21)    <= sub_wire15(21);
	sub_wire2(18, 22)    <= sub_wire15(22);
	sub_wire2(18, 23)    <= sub_wire15(23);
	sub_wire2(18, 24)    <= sub_wire15(24);
	sub_wire2(18, 25)    <= sub_wire15(25);
	sub_wire2(18, 26)    <= sub_wire15(26);
	sub_wire2(18, 27)    <= sub_wire15(27);
	sub_wire2(18, 28)    <= sub_wire15(28);
	sub_wire2(18, 29)    <= sub_wire15(29);
	sub_wire2(18, 30)    <= sub_wire15(30);
	sub_wire2(18, 31)    <= sub_wire15(31);
	sub_wire2(17, 0)    <= sub_wire16(0);
	sub_wire2(17, 1)    <= sub_wire16(1);
	sub_wire2(17, 2)    <= sub_wire16(2);
	sub_wire2(17, 3)    <= sub_wire16(3);
	sub_wire2(17, 4)    <= sub_wire16(4);
	sub_wire2(17, 5)    <= sub_wire16(5);
	sub_wire2(17, 6)    <= sub_wire16(6);
	sub_wire2(17, 7)    <= sub_wire16(7);
	sub_wire2(17, 8)    <= sub_wire16(8);
	sub_wire2(17, 9)    <= sub_wire16(9);
	sub_wire2(17, 10)    <= sub_wire16(10);
	sub_wire2(17, 11)    <= sub_wire16(11);
	sub_wire2(17, 12)    <= sub_wire16(12);
	sub_wire2(17, 13)    <= sub_wire16(13);
	sub_wire2(17, 14)    <= sub_wire16(14);
	sub_wire2(17, 15)    <= sub_wire16(15);
	sub_wire2(17, 16)    <= sub_wire16(16);
	sub_wire2(17, 17)    <= sub_wire16(17);
	sub_wire2(17, 18)    <= sub_wire16(18);
	sub_wire2(17, 19)    <= sub_wire16(19);
	sub_wire2(17, 20)    <= sub_wire16(20);
	sub_wire2(17, 21)    <= sub_wire16(21);
	sub_wire2(17, 22)    <= sub_wire16(22);
	sub_wire2(17, 23)    <= sub_wire16(23);
	sub_wire2(17, 24)    <= sub_wire16(24);
	sub_wire2(17, 25)    <= sub_wire16(25);
	sub_wire2(17, 26)    <= sub_wire16(26);
	sub_wire2(17, 27)    <= sub_wire16(27);
	sub_wire2(17, 28)    <= sub_wire16(28);
	sub_wire2(17, 29)    <= sub_wire16(29);
	sub_wire2(17, 30)    <= sub_wire16(30);
	sub_wire2(17, 31)    <= sub_wire16(31);
	sub_wire2(16, 0)    <= sub_wire17(0);
	sub_wire2(16, 1)    <= sub_wire17(1);
	sub_wire2(16, 2)    <= sub_wire17(2);
	sub_wire2(16, 3)    <= sub_wire17(3);
	sub_wire2(16, 4)    <= sub_wire17(4);
	sub_wire2(16, 5)    <= sub_wire17(5);
	sub_wire2(16, 6)    <= sub_wire17(6);
	sub_wire2(16, 7)    <= sub_wire17(7);
	sub_wire2(16, 8)    <= sub_wire17(8);
	sub_wire2(16, 9)    <= sub_wire17(9);
	sub_wire2(16, 10)    <= sub_wire17(10);
	sub_wire2(16, 11)    <= sub_wire17(11);
	sub_wire2(16, 12)    <= sub_wire17(12);
	sub_wire2(16, 13)    <= sub_wire17(13);
	sub_wire2(16, 14)    <= sub_wire17(14);
	sub_wire2(16, 15)    <= sub_wire17(15);
	sub_wire2(16, 16)    <= sub_wire17(16);
	sub_wire2(16, 17)    <= sub_wire17(17);
	sub_wire2(16, 18)    <= sub_wire17(18);
	sub_wire2(16, 19)    <= sub_wire17(19);
	sub_wire2(16, 20)    <= sub_wire17(20);
	sub_wire2(16, 21)    <= sub_wire17(21);
	sub_wire2(16, 22)    <= sub_wire17(22);
	sub_wire2(16, 23)    <= sub_wire17(23);
	sub_wire2(16, 24)    <= sub_wire17(24);
	sub_wire2(16, 25)    <= sub_wire17(25);
	sub_wire2(16, 26)    <= sub_wire17(26);
	sub_wire2(16, 27)    <= sub_wire17(27);
	sub_wire2(16, 28)    <= sub_wire17(28);
	sub_wire2(16, 29)    <= sub_wire17(29);
	sub_wire2(16, 30)    <= sub_wire17(30);
	sub_wire2(16, 31)    <= sub_wire17(31);
	sub_wire2(15, 0)    <= sub_wire18(0);
	sub_wire2(15, 1)    <= sub_wire18(1);
	sub_wire2(15, 2)    <= sub_wire18(2);
	sub_wire2(15, 3)    <= sub_wire18(3);
	sub_wire2(15, 4)    <= sub_wire18(4);
	sub_wire2(15, 5)    <= sub_wire18(5);
	sub_wire2(15, 6)    <= sub_wire18(6);
	sub_wire2(15, 7)    <= sub_wire18(7);
	sub_wire2(15, 8)    <= sub_wire18(8);
	sub_wire2(15, 9)    <= sub_wire18(9);
	sub_wire2(15, 10)    <= sub_wire18(10);
	sub_wire2(15, 11)    <= sub_wire18(11);
	sub_wire2(15, 12)    <= sub_wire18(12);
	sub_wire2(15, 13)    <= sub_wire18(13);
	sub_wire2(15, 14)    <= sub_wire18(14);
	sub_wire2(15, 15)    <= sub_wire18(15);
	sub_wire2(15, 16)    <= sub_wire18(16);
	sub_wire2(15, 17)    <= sub_wire18(17);
	sub_wire2(15, 18)    <= sub_wire18(18);
	sub_wire2(15, 19)    <= sub_wire18(19);
	sub_wire2(15, 20)    <= sub_wire18(20);
	sub_wire2(15, 21)    <= sub_wire18(21);
	sub_wire2(15, 22)    <= sub_wire18(22);
	sub_wire2(15, 23)    <= sub_wire18(23);
	sub_wire2(15, 24)    <= sub_wire18(24);
	sub_wire2(15, 25)    <= sub_wire18(25);
	sub_wire2(15, 26)    <= sub_wire18(26);
	sub_wire2(15, 27)    <= sub_wire18(27);
	sub_wire2(15, 28)    <= sub_wire18(28);
	sub_wire2(15, 29)    <= sub_wire18(29);
	sub_wire2(15, 30)    <= sub_wire18(30);
	sub_wire2(15, 31)    <= sub_wire18(31);
	sub_wire2(14, 0)    <= sub_wire19(0);
	sub_wire2(14, 1)    <= sub_wire19(1);
	sub_wire2(14, 2)    <= sub_wire19(2);
	sub_wire2(14, 3)    <= sub_wire19(3);
	sub_wire2(14, 4)    <= sub_wire19(4);
	sub_wire2(14, 5)    <= sub_wire19(5);
	sub_wire2(14, 6)    <= sub_wire19(6);
	sub_wire2(14, 7)    <= sub_wire19(7);
	sub_wire2(14, 8)    <= sub_wire19(8);
	sub_wire2(14, 9)    <= sub_wire19(9);
	sub_wire2(14, 10)    <= sub_wire19(10);
	sub_wire2(14, 11)    <= sub_wire19(11);
	sub_wire2(14, 12)    <= sub_wire19(12);
	sub_wire2(14, 13)    <= sub_wire19(13);
	sub_wire2(14, 14)    <= sub_wire19(14);
	sub_wire2(14, 15)    <= sub_wire19(15);
	sub_wire2(14, 16)    <= sub_wire19(16);
	sub_wire2(14, 17)    <= sub_wire19(17);
	sub_wire2(14, 18)    <= sub_wire19(18);
	sub_wire2(14, 19)    <= sub_wire19(19);
	sub_wire2(14, 20)    <= sub_wire19(20);
	sub_wire2(14, 21)    <= sub_wire19(21);
	sub_wire2(14, 22)    <= sub_wire19(22);
	sub_wire2(14, 23)    <= sub_wire19(23);
	sub_wire2(14, 24)    <= sub_wire19(24);
	sub_wire2(14, 25)    <= sub_wire19(25);
	sub_wire2(14, 26)    <= sub_wire19(26);
	sub_wire2(14, 27)    <= sub_wire19(27);
	sub_wire2(14, 28)    <= sub_wire19(28);
	sub_wire2(14, 29)    <= sub_wire19(29);
	sub_wire2(14, 30)    <= sub_wire19(30);
	sub_wire2(14, 31)    <= sub_wire19(31);
	sub_wire2(13, 0)    <= sub_wire20(0);
	sub_wire2(13, 1)    <= sub_wire20(1);
	sub_wire2(13, 2)    <= sub_wire20(2);
	sub_wire2(13, 3)    <= sub_wire20(3);
	sub_wire2(13, 4)    <= sub_wire20(4);
	sub_wire2(13, 5)    <= sub_wire20(5);
	sub_wire2(13, 6)    <= sub_wire20(6);
	sub_wire2(13, 7)    <= sub_wire20(7);
	sub_wire2(13, 8)    <= sub_wire20(8);
	sub_wire2(13, 9)    <= sub_wire20(9);
	sub_wire2(13, 10)    <= sub_wire20(10);
	sub_wire2(13, 11)    <= sub_wire20(11);
	sub_wire2(13, 12)    <= sub_wire20(12);
	sub_wire2(13, 13)    <= sub_wire20(13);
	sub_wire2(13, 14)    <= sub_wire20(14);
	sub_wire2(13, 15)    <= sub_wire20(15);
	sub_wire2(13, 16)    <= sub_wire20(16);
	sub_wire2(13, 17)    <= sub_wire20(17);
	sub_wire2(13, 18)    <= sub_wire20(18);
	sub_wire2(13, 19)    <= sub_wire20(19);
	sub_wire2(13, 20)    <= sub_wire20(20);
	sub_wire2(13, 21)    <= sub_wire20(21);
	sub_wire2(13, 22)    <= sub_wire20(22);
	sub_wire2(13, 23)    <= sub_wire20(23);
	sub_wire2(13, 24)    <= sub_wire20(24);
	sub_wire2(13, 25)    <= sub_wire20(25);
	sub_wire2(13, 26)    <= sub_wire20(26);
	sub_wire2(13, 27)    <= sub_wire20(27);
	sub_wire2(13, 28)    <= sub_wire20(28);
	sub_wire2(13, 29)    <= sub_wire20(29);
	sub_wire2(13, 30)    <= sub_wire20(30);
	sub_wire2(13, 31)    <= sub_wire20(31);
	sub_wire2(12, 0)    <= sub_wire21(0);
	sub_wire2(12, 1)    <= sub_wire21(1);
	sub_wire2(12, 2)    <= sub_wire21(2);
	sub_wire2(12, 3)    <= sub_wire21(3);
	sub_wire2(12, 4)    <= sub_wire21(4);
	sub_wire2(12, 5)    <= sub_wire21(5);
	sub_wire2(12, 6)    <= sub_wire21(6);
	sub_wire2(12, 7)    <= sub_wire21(7);
	sub_wire2(12, 8)    <= sub_wire21(8);
	sub_wire2(12, 9)    <= sub_wire21(9);
	sub_wire2(12, 10)    <= sub_wire21(10);
	sub_wire2(12, 11)    <= sub_wire21(11);
	sub_wire2(12, 12)    <= sub_wire21(12);
	sub_wire2(12, 13)    <= sub_wire21(13);
	sub_wire2(12, 14)    <= sub_wire21(14);
	sub_wire2(12, 15)    <= sub_wire21(15);
	sub_wire2(12, 16)    <= sub_wire21(16);
	sub_wire2(12, 17)    <= sub_wire21(17);
	sub_wire2(12, 18)    <= sub_wire21(18);
	sub_wire2(12, 19)    <= sub_wire21(19);
	sub_wire2(12, 20)    <= sub_wire21(20);
	sub_wire2(12, 21)    <= sub_wire21(21);
	sub_wire2(12, 22)    <= sub_wire21(22);
	sub_wire2(12, 23)    <= sub_wire21(23);
	sub_wire2(12, 24)    <= sub_wire21(24);
	sub_wire2(12, 25)    <= sub_wire21(25);
	sub_wire2(12, 26)    <= sub_wire21(26);
	sub_wire2(12, 27)    <= sub_wire21(27);
	sub_wire2(12, 28)    <= sub_wire21(28);
	sub_wire2(12, 29)    <= sub_wire21(29);
	sub_wire2(12, 30)    <= sub_wire21(30);
	sub_wire2(12, 31)    <= sub_wire21(31);
	sub_wire2(11, 0)    <= sub_wire22(0);
	sub_wire2(11, 1)    <= sub_wire22(1);
	sub_wire2(11, 2)    <= sub_wire22(2);
	sub_wire2(11, 3)    <= sub_wire22(3);
	sub_wire2(11, 4)    <= sub_wire22(4);
	sub_wire2(11, 5)    <= sub_wire22(5);
	sub_wire2(11, 6)    <= sub_wire22(6);
	sub_wire2(11, 7)    <= sub_wire22(7);
	sub_wire2(11, 8)    <= sub_wire22(8);
	sub_wire2(11, 9)    <= sub_wire22(9);
	sub_wire2(11, 10)    <= sub_wire22(10);
	sub_wire2(11, 11)    <= sub_wire22(11);
	sub_wire2(11, 12)    <= sub_wire22(12);
	sub_wire2(11, 13)    <= sub_wire22(13);
	sub_wire2(11, 14)    <= sub_wire22(14);
	sub_wire2(11, 15)    <= sub_wire22(15);
	sub_wire2(11, 16)    <= sub_wire22(16);
	sub_wire2(11, 17)    <= sub_wire22(17);
	sub_wire2(11, 18)    <= sub_wire22(18);
	sub_wire2(11, 19)    <= sub_wire22(19);
	sub_wire2(11, 20)    <= sub_wire22(20);
	sub_wire2(11, 21)    <= sub_wire22(21);
	sub_wire2(11, 22)    <= sub_wire22(22);
	sub_wire2(11, 23)    <= sub_wire22(23);
	sub_wire2(11, 24)    <= sub_wire22(24);
	sub_wire2(11, 25)    <= sub_wire22(25);
	sub_wire2(11, 26)    <= sub_wire22(26);
	sub_wire2(11, 27)    <= sub_wire22(27);
	sub_wire2(11, 28)    <= sub_wire22(28);
	sub_wire2(11, 29)    <= sub_wire22(29);
	sub_wire2(11, 30)    <= sub_wire22(30);
	sub_wire2(11, 31)    <= sub_wire22(31);
	sub_wire2(10, 0)    <= sub_wire23(0);
	sub_wire2(10, 1)    <= sub_wire23(1);
	sub_wire2(10, 2)    <= sub_wire23(2);
	sub_wire2(10, 3)    <= sub_wire23(3);
	sub_wire2(10, 4)    <= sub_wire23(4);
	sub_wire2(10, 5)    <= sub_wire23(5);
	sub_wire2(10, 6)    <= sub_wire23(6);
	sub_wire2(10, 7)    <= sub_wire23(7);
	sub_wire2(10, 8)    <= sub_wire23(8);
	sub_wire2(10, 9)    <= sub_wire23(9);
	sub_wire2(10, 10)    <= sub_wire23(10);
	sub_wire2(10, 11)    <= sub_wire23(11);
	sub_wire2(10, 12)    <= sub_wire23(12);
	sub_wire2(10, 13)    <= sub_wire23(13);
	sub_wire2(10, 14)    <= sub_wire23(14);
	sub_wire2(10, 15)    <= sub_wire23(15);
	sub_wire2(10, 16)    <= sub_wire23(16);
	sub_wire2(10, 17)    <= sub_wire23(17);
	sub_wire2(10, 18)    <= sub_wire23(18);
	sub_wire2(10, 19)    <= sub_wire23(19);
	sub_wire2(10, 20)    <= sub_wire23(20);
	sub_wire2(10, 21)    <= sub_wire23(21);
	sub_wire2(10, 22)    <= sub_wire23(22);
	sub_wire2(10, 23)    <= sub_wire23(23);
	sub_wire2(10, 24)    <= sub_wire23(24);
	sub_wire2(10, 25)    <= sub_wire23(25);
	sub_wire2(10, 26)    <= sub_wire23(26);
	sub_wire2(10, 27)    <= sub_wire23(27);
	sub_wire2(10, 28)    <= sub_wire23(28);
	sub_wire2(10, 29)    <= sub_wire23(29);
	sub_wire2(10, 30)    <= sub_wire23(30);
	sub_wire2(10, 31)    <= sub_wire23(31);
	sub_wire2(9, 0)    <= sub_wire24(0);
	sub_wire2(9, 1)    <= sub_wire24(1);
	sub_wire2(9, 2)    <= sub_wire24(2);
	sub_wire2(9, 3)    <= sub_wire24(3);
	sub_wire2(9, 4)    <= sub_wire24(4);
	sub_wire2(9, 5)    <= sub_wire24(5);
	sub_wire2(9, 6)    <= sub_wire24(6);
	sub_wire2(9, 7)    <= sub_wire24(7);
	sub_wire2(9, 8)    <= sub_wire24(8);
	sub_wire2(9, 9)    <= sub_wire24(9);
	sub_wire2(9, 10)    <= sub_wire24(10);
	sub_wire2(9, 11)    <= sub_wire24(11);
	sub_wire2(9, 12)    <= sub_wire24(12);
	sub_wire2(9, 13)    <= sub_wire24(13);
	sub_wire2(9, 14)    <= sub_wire24(14);
	sub_wire2(9, 15)    <= sub_wire24(15);
	sub_wire2(9, 16)    <= sub_wire24(16);
	sub_wire2(9, 17)    <= sub_wire24(17);
	sub_wire2(9, 18)    <= sub_wire24(18);
	sub_wire2(9, 19)    <= sub_wire24(19);
	sub_wire2(9, 20)    <= sub_wire24(20);
	sub_wire2(9, 21)    <= sub_wire24(21);
	sub_wire2(9, 22)    <= sub_wire24(22);
	sub_wire2(9, 23)    <= sub_wire24(23);
	sub_wire2(9, 24)    <= sub_wire24(24);
	sub_wire2(9, 25)    <= sub_wire24(25);
	sub_wire2(9, 26)    <= sub_wire24(26);
	sub_wire2(9, 27)    <= sub_wire24(27);
	sub_wire2(9, 28)    <= sub_wire24(28);
	sub_wire2(9, 29)    <= sub_wire24(29);
	sub_wire2(9, 30)    <= sub_wire24(30);
	sub_wire2(9, 31)    <= sub_wire24(31);
	sub_wire2(8, 0)    <= sub_wire25(0);
	sub_wire2(8, 1)    <= sub_wire25(1);
	sub_wire2(8, 2)    <= sub_wire25(2);
	sub_wire2(8, 3)    <= sub_wire25(3);
	sub_wire2(8, 4)    <= sub_wire25(4);
	sub_wire2(8, 5)    <= sub_wire25(5);
	sub_wire2(8, 6)    <= sub_wire25(6);
	sub_wire2(8, 7)    <= sub_wire25(7);
	sub_wire2(8, 8)    <= sub_wire25(8);
	sub_wire2(8, 9)    <= sub_wire25(9);
	sub_wire2(8, 10)    <= sub_wire25(10);
	sub_wire2(8, 11)    <= sub_wire25(11);
	sub_wire2(8, 12)    <= sub_wire25(12);
	sub_wire2(8, 13)    <= sub_wire25(13);
	sub_wire2(8, 14)    <= sub_wire25(14);
	sub_wire2(8, 15)    <= sub_wire25(15);
	sub_wire2(8, 16)    <= sub_wire25(16);
	sub_wire2(8, 17)    <= sub_wire25(17);
	sub_wire2(8, 18)    <= sub_wire25(18);
	sub_wire2(8, 19)    <= sub_wire25(19);
	sub_wire2(8, 20)    <= sub_wire25(20);
	sub_wire2(8, 21)    <= sub_wire25(21);
	sub_wire2(8, 22)    <= sub_wire25(22);
	sub_wire2(8, 23)    <= sub_wire25(23);
	sub_wire2(8, 24)    <= sub_wire25(24);
	sub_wire2(8, 25)    <= sub_wire25(25);
	sub_wire2(8, 26)    <= sub_wire25(26);
	sub_wire2(8, 27)    <= sub_wire25(27);
	sub_wire2(8, 28)    <= sub_wire25(28);
	sub_wire2(8, 29)    <= sub_wire25(29);
	sub_wire2(8, 30)    <= sub_wire25(30);
	sub_wire2(8, 31)    <= sub_wire25(31);
	sub_wire2(7, 0)    <= sub_wire26(0);
	sub_wire2(7, 1)    <= sub_wire26(1);
	sub_wire2(7, 2)    <= sub_wire26(2);
	sub_wire2(7, 3)    <= sub_wire26(3);
	sub_wire2(7, 4)    <= sub_wire26(4);
	sub_wire2(7, 5)    <= sub_wire26(5);
	sub_wire2(7, 6)    <= sub_wire26(6);
	sub_wire2(7, 7)    <= sub_wire26(7);
	sub_wire2(7, 8)    <= sub_wire26(8);
	sub_wire2(7, 9)    <= sub_wire26(9);
	sub_wire2(7, 10)    <= sub_wire26(10);
	sub_wire2(7, 11)    <= sub_wire26(11);
	sub_wire2(7, 12)    <= sub_wire26(12);
	sub_wire2(7, 13)    <= sub_wire26(13);
	sub_wire2(7, 14)    <= sub_wire26(14);
	sub_wire2(7, 15)    <= sub_wire26(15);
	sub_wire2(7, 16)    <= sub_wire26(16);
	sub_wire2(7, 17)    <= sub_wire26(17);
	sub_wire2(7, 18)    <= sub_wire26(18);
	sub_wire2(7, 19)    <= sub_wire26(19);
	sub_wire2(7, 20)    <= sub_wire26(20);
	sub_wire2(7, 21)    <= sub_wire26(21);
	sub_wire2(7, 22)    <= sub_wire26(22);
	sub_wire2(7, 23)    <= sub_wire26(23);
	sub_wire2(7, 24)    <= sub_wire26(24);
	sub_wire2(7, 25)    <= sub_wire26(25);
	sub_wire2(7, 26)    <= sub_wire26(26);
	sub_wire2(7, 27)    <= sub_wire26(27);
	sub_wire2(7, 28)    <= sub_wire26(28);
	sub_wire2(7, 29)    <= sub_wire26(29);
	sub_wire2(7, 30)    <= sub_wire26(30);
	sub_wire2(7, 31)    <= sub_wire26(31);
	sub_wire2(6, 0)    <= sub_wire27(0);
	sub_wire2(6, 1)    <= sub_wire27(1);
	sub_wire2(6, 2)    <= sub_wire27(2);
	sub_wire2(6, 3)    <= sub_wire27(3);
	sub_wire2(6, 4)    <= sub_wire27(4);
	sub_wire2(6, 5)    <= sub_wire27(5);
	sub_wire2(6, 6)    <= sub_wire27(6);
	sub_wire2(6, 7)    <= sub_wire27(7);
	sub_wire2(6, 8)    <= sub_wire27(8);
	sub_wire2(6, 9)    <= sub_wire27(9);
	sub_wire2(6, 10)    <= sub_wire27(10);
	sub_wire2(6, 11)    <= sub_wire27(11);
	sub_wire2(6, 12)    <= sub_wire27(12);
	sub_wire2(6, 13)    <= sub_wire27(13);
	sub_wire2(6, 14)    <= sub_wire27(14);
	sub_wire2(6, 15)    <= sub_wire27(15);
	sub_wire2(6, 16)    <= sub_wire27(16);
	sub_wire2(6, 17)    <= sub_wire27(17);
	sub_wire2(6, 18)    <= sub_wire27(18);
	sub_wire2(6, 19)    <= sub_wire27(19);
	sub_wire2(6, 20)    <= sub_wire27(20);
	sub_wire2(6, 21)    <= sub_wire27(21);
	sub_wire2(6, 22)    <= sub_wire27(22);
	sub_wire2(6, 23)    <= sub_wire27(23);
	sub_wire2(6, 24)    <= sub_wire27(24);
	sub_wire2(6, 25)    <= sub_wire27(25);
	sub_wire2(6, 26)    <= sub_wire27(26);
	sub_wire2(6, 27)    <= sub_wire27(27);
	sub_wire2(6, 28)    <= sub_wire27(28);
	sub_wire2(6, 29)    <= sub_wire27(29);
	sub_wire2(6, 30)    <= sub_wire27(30);
	sub_wire2(6, 31)    <= sub_wire27(31);
	sub_wire2(5, 0)    <= sub_wire28(0);
	sub_wire2(5, 1)    <= sub_wire28(1);
	sub_wire2(5, 2)    <= sub_wire28(2);
	sub_wire2(5, 3)    <= sub_wire28(3);
	sub_wire2(5, 4)    <= sub_wire28(4);
	sub_wire2(5, 5)    <= sub_wire28(5);
	sub_wire2(5, 6)    <= sub_wire28(6);
	sub_wire2(5, 7)    <= sub_wire28(7);
	sub_wire2(5, 8)    <= sub_wire28(8);
	sub_wire2(5, 9)    <= sub_wire28(9);
	sub_wire2(5, 10)    <= sub_wire28(10);
	sub_wire2(5, 11)    <= sub_wire28(11);
	sub_wire2(5, 12)    <= sub_wire28(12);
	sub_wire2(5, 13)    <= sub_wire28(13);
	sub_wire2(5, 14)    <= sub_wire28(14);
	sub_wire2(5, 15)    <= sub_wire28(15);
	sub_wire2(5, 16)    <= sub_wire28(16);
	sub_wire2(5, 17)    <= sub_wire28(17);
	sub_wire2(5, 18)    <= sub_wire28(18);
	sub_wire2(5, 19)    <= sub_wire28(19);
	sub_wire2(5, 20)    <= sub_wire28(20);
	sub_wire2(5, 21)    <= sub_wire28(21);
	sub_wire2(5, 22)    <= sub_wire28(22);
	sub_wire2(5, 23)    <= sub_wire28(23);
	sub_wire2(5, 24)    <= sub_wire28(24);
	sub_wire2(5, 25)    <= sub_wire28(25);
	sub_wire2(5, 26)    <= sub_wire28(26);
	sub_wire2(5, 27)    <= sub_wire28(27);
	sub_wire2(5, 28)    <= sub_wire28(28);
	sub_wire2(5, 29)    <= sub_wire28(29);
	sub_wire2(5, 30)    <= sub_wire28(30);
	sub_wire2(5, 31)    <= sub_wire28(31);
	sub_wire2(4, 0)    <= sub_wire29(0);
	sub_wire2(4, 1)    <= sub_wire29(1);
	sub_wire2(4, 2)    <= sub_wire29(2);
	sub_wire2(4, 3)    <= sub_wire29(3);
	sub_wire2(4, 4)    <= sub_wire29(4);
	sub_wire2(4, 5)    <= sub_wire29(5);
	sub_wire2(4, 6)    <= sub_wire29(6);
	sub_wire2(4, 7)    <= sub_wire29(7);
	sub_wire2(4, 8)    <= sub_wire29(8);
	sub_wire2(4, 9)    <= sub_wire29(9);
	sub_wire2(4, 10)    <= sub_wire29(10);
	sub_wire2(4, 11)    <= sub_wire29(11);
	sub_wire2(4, 12)    <= sub_wire29(12);
	sub_wire2(4, 13)    <= sub_wire29(13);
	sub_wire2(4, 14)    <= sub_wire29(14);
	sub_wire2(4, 15)    <= sub_wire29(15);
	sub_wire2(4, 16)    <= sub_wire29(16);
	sub_wire2(4, 17)    <= sub_wire29(17);
	sub_wire2(4, 18)    <= sub_wire29(18);
	sub_wire2(4, 19)    <= sub_wire29(19);
	sub_wire2(4, 20)    <= sub_wire29(20);
	sub_wire2(4, 21)    <= sub_wire29(21);
	sub_wire2(4, 22)    <= sub_wire29(22);
	sub_wire2(4, 23)    <= sub_wire29(23);
	sub_wire2(4, 24)    <= sub_wire29(24);
	sub_wire2(4, 25)    <= sub_wire29(25);
	sub_wire2(4, 26)    <= sub_wire29(26);
	sub_wire2(4, 27)    <= sub_wire29(27);
	sub_wire2(4, 28)    <= sub_wire29(28);
	sub_wire2(4, 29)    <= sub_wire29(29);
	sub_wire2(4, 30)    <= sub_wire29(30);
	sub_wire2(4, 31)    <= sub_wire29(31);
	sub_wire2(3, 0)    <= sub_wire30(0);
	sub_wire2(3, 1)    <= sub_wire30(1);
	sub_wire2(3, 2)    <= sub_wire30(2);
	sub_wire2(3, 3)    <= sub_wire30(3);
	sub_wire2(3, 4)    <= sub_wire30(4);
	sub_wire2(3, 5)    <= sub_wire30(5);
	sub_wire2(3, 6)    <= sub_wire30(6);
	sub_wire2(3, 7)    <= sub_wire30(7);
	sub_wire2(3, 8)    <= sub_wire30(8);
	sub_wire2(3, 9)    <= sub_wire30(9);
	sub_wire2(3, 10)    <= sub_wire30(10);
	sub_wire2(3, 11)    <= sub_wire30(11);
	sub_wire2(3, 12)    <= sub_wire30(12);
	sub_wire2(3, 13)    <= sub_wire30(13);
	sub_wire2(3, 14)    <= sub_wire30(14);
	sub_wire2(3, 15)    <= sub_wire30(15);
	sub_wire2(3, 16)    <= sub_wire30(16);
	sub_wire2(3, 17)    <= sub_wire30(17);
	sub_wire2(3, 18)    <= sub_wire30(18);
	sub_wire2(3, 19)    <= sub_wire30(19);
	sub_wire2(3, 20)    <= sub_wire30(20);
	sub_wire2(3, 21)    <= sub_wire30(21);
	sub_wire2(3, 22)    <= sub_wire30(22);
	sub_wire2(3, 23)    <= sub_wire30(23);
	sub_wire2(3, 24)    <= sub_wire30(24);
	sub_wire2(3, 25)    <= sub_wire30(25);
	sub_wire2(3, 26)    <= sub_wire30(26);
	sub_wire2(3, 27)    <= sub_wire30(27);
	sub_wire2(3, 28)    <= sub_wire30(28);
	sub_wire2(3, 29)    <= sub_wire30(29);
	sub_wire2(3, 30)    <= sub_wire30(30);
	sub_wire2(3, 31)    <= sub_wire30(31);
	sub_wire2(2, 0)    <= sub_wire31(0);
	sub_wire2(2, 1)    <= sub_wire31(1);
	sub_wire2(2, 2)    <= sub_wire31(2);
	sub_wire2(2, 3)    <= sub_wire31(3);
	sub_wire2(2, 4)    <= sub_wire31(4);
	sub_wire2(2, 5)    <= sub_wire31(5);
	sub_wire2(2, 6)    <= sub_wire31(6);
	sub_wire2(2, 7)    <= sub_wire31(7);
	sub_wire2(2, 8)    <= sub_wire31(8);
	sub_wire2(2, 9)    <= sub_wire31(9);
	sub_wire2(2, 10)    <= sub_wire31(10);
	sub_wire2(2, 11)    <= sub_wire31(11);
	sub_wire2(2, 12)    <= sub_wire31(12);
	sub_wire2(2, 13)    <= sub_wire31(13);
	sub_wire2(2, 14)    <= sub_wire31(14);
	sub_wire2(2, 15)    <= sub_wire31(15);
	sub_wire2(2, 16)    <= sub_wire31(16);
	sub_wire2(2, 17)    <= sub_wire31(17);
	sub_wire2(2, 18)    <= sub_wire31(18);
	sub_wire2(2, 19)    <= sub_wire31(19);
	sub_wire2(2, 20)    <= sub_wire31(20);
	sub_wire2(2, 21)    <= sub_wire31(21);
	sub_wire2(2, 22)    <= sub_wire31(22);
	sub_wire2(2, 23)    <= sub_wire31(23);
	sub_wire2(2, 24)    <= sub_wire31(24);
	sub_wire2(2, 25)    <= sub_wire31(25);
	sub_wire2(2, 26)    <= sub_wire31(26);
	sub_wire2(2, 27)    <= sub_wire31(27);
	sub_wire2(2, 28)    <= sub_wire31(28);
	sub_wire2(2, 29)    <= sub_wire31(29);
	sub_wire2(2, 30)    <= sub_wire31(30);
	sub_wire2(2, 31)    <= sub_wire31(31);
	sub_wire2(1, 0)    <= sub_wire32(0);
	sub_wire2(1, 1)    <= sub_wire32(1);
	sub_wire2(1, 2)    <= sub_wire32(2);
	sub_wire2(1, 3)    <= sub_wire32(3);
	sub_wire2(1, 4)    <= sub_wire32(4);
	sub_wire2(1, 5)    <= sub_wire32(5);
	sub_wire2(1, 6)    <= sub_wire32(6);
	sub_wire2(1, 7)    <= sub_wire32(7);
	sub_wire2(1, 8)    <= sub_wire32(8);
	sub_wire2(1, 9)    <= sub_wire32(9);
	sub_wire2(1, 10)    <= sub_wire32(10);
	sub_wire2(1, 11)    <= sub_wire32(11);
	sub_wire2(1, 12)    <= sub_wire32(12);
	sub_wire2(1, 13)    <= sub_wire32(13);
	sub_wire2(1, 14)    <= sub_wire32(14);
	sub_wire2(1, 15)    <= sub_wire32(15);
	sub_wire2(1, 16)    <= sub_wire32(16);
	sub_wire2(1, 17)    <= sub_wire32(17);
	sub_wire2(1, 18)    <= sub_wire32(18);
	sub_wire2(1, 19)    <= sub_wire32(19);
	sub_wire2(1, 20)    <= sub_wire32(20);
	sub_wire2(1, 21)    <= sub_wire32(21);
	sub_wire2(1, 22)    <= sub_wire32(22);
	sub_wire2(1, 23)    <= sub_wire32(23);
	sub_wire2(1, 24)    <= sub_wire32(24);
	sub_wire2(1, 25)    <= sub_wire32(25);
	sub_wire2(1, 26)    <= sub_wire32(26);
	sub_wire2(1, 27)    <= sub_wire32(27);
	sub_wire2(1, 28)    <= sub_wire32(28);
	sub_wire2(1, 29)    <= sub_wire32(29);
	sub_wire2(1, 30)    <= sub_wire32(30);
	sub_wire2(1, 31)    <= sub_wire32(31);
	sub_wire2(0, 0)    <= sub_wire33(0);
	sub_wire2(0, 1)    <= sub_wire33(1);
	sub_wire2(0, 2)    <= sub_wire33(2);
	sub_wire2(0, 3)    <= sub_wire33(3);
	sub_wire2(0, 4)    <= sub_wire33(4);
	sub_wire2(0, 5)    <= sub_wire33(5);
	sub_wire2(0, 6)    <= sub_wire33(6);
	sub_wire2(0, 7)    <= sub_wire33(7);
	sub_wire2(0, 8)    <= sub_wire33(8);
	sub_wire2(0, 9)    <= sub_wire33(9);
	sub_wire2(0, 10)    <= sub_wire33(10);
	sub_wire2(0, 11)    <= sub_wire33(11);
	sub_wire2(0, 12)    <= sub_wire33(12);
	sub_wire2(0, 13)    <= sub_wire33(13);
	sub_wire2(0, 14)    <= sub_wire33(14);
	sub_wire2(0, 15)    <= sub_wire33(15);
	sub_wire2(0, 16)    <= sub_wire33(16);
	sub_wire2(0, 17)    <= sub_wire33(17);
	sub_wire2(0, 18)    <= sub_wire33(18);
	sub_wire2(0, 19)    <= sub_wire33(19);
	sub_wire2(0, 20)    <= sub_wire33(20);
	sub_wire2(0, 21)    <= sub_wire33(21);
	sub_wire2(0, 22)    <= sub_wire33(22);
	sub_wire2(0, 23)    <= sub_wire33(23);
	sub_wire2(0, 24)    <= sub_wire33(24);
	sub_wire2(0, 25)    <= sub_wire33(25);
	sub_wire2(0, 26)    <= sub_wire33(26);
	sub_wire2(0, 27)    <= sub_wire33(27);
	sub_wire2(0, 28)    <= sub_wire33(28);
	sub_wire2(0, 29)    <= sub_wire33(29);
	sub_wire2(0, 30)    <= sub_wire33(30);
	sub_wire2(0, 31)    <= sub_wire33(31);

	LPM_MUX_component : LPM_MUX
	GENERIC MAP (
		lpm_size => 32,
		lpm_type => "LPM_MUX",
		lpm_width => 32,
		lpm_widths => 5
	)
	PORT MAP (
		data => sub_wire2,
		sel => sel,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "5"
-- Retrieval info: USED_PORT: data0x 0 0 32 0 INPUT NODEFVAL "data0x[31..0]"
-- Retrieval info: USED_PORT: data10x 0 0 32 0 INPUT NODEFVAL "data10x[31..0]"
-- Retrieval info: USED_PORT: data11x 0 0 32 0 INPUT NODEFVAL "data11x[31..0]"
-- Retrieval info: USED_PORT: data12x 0 0 32 0 INPUT NODEFVAL "data12x[31..0]"
-- Retrieval info: USED_PORT: data13x 0 0 32 0 INPUT NODEFVAL "data13x[31..0]"
-- Retrieval info: USED_PORT: data14x 0 0 32 0 INPUT NODEFVAL "data14x[31..0]"
-- Retrieval info: USED_PORT: data15x 0 0 32 0 INPUT NODEFVAL "data15x[31..0]"
-- Retrieval info: USED_PORT: data16x 0 0 32 0 INPUT NODEFVAL "data16x[31..0]"
-- Retrieval info: USED_PORT: data17x 0 0 32 0 INPUT NODEFVAL "data17x[31..0]"
-- Retrieval info: USED_PORT: data18x 0 0 32 0 INPUT NODEFVAL "data18x[31..0]"
-- Retrieval info: USED_PORT: data19x 0 0 32 0 INPUT NODEFVAL "data19x[31..0]"
-- Retrieval info: USED_PORT: data1x 0 0 32 0 INPUT NODEFVAL "data1x[31..0]"
-- Retrieval info: USED_PORT: data20x 0 0 32 0 INPUT NODEFVAL "data20x[31..0]"
-- Retrieval info: USED_PORT: data21x 0 0 32 0 INPUT NODEFVAL "data21x[31..0]"
-- Retrieval info: USED_PORT: data22x 0 0 32 0 INPUT NODEFVAL "data22x[31..0]"
-- Retrieval info: USED_PORT: data23x 0 0 32 0 INPUT NODEFVAL "data23x[31..0]"
-- Retrieval info: USED_PORT: data24x 0 0 32 0 INPUT NODEFVAL "data24x[31..0]"
-- Retrieval info: USED_PORT: data25x 0 0 32 0 INPUT NODEFVAL "data25x[31..0]"
-- Retrieval info: USED_PORT: data26x 0 0 32 0 INPUT NODEFVAL "data26x[31..0]"
-- Retrieval info: USED_PORT: data27x 0 0 32 0 INPUT NODEFVAL "data27x[31..0]"
-- Retrieval info: USED_PORT: data28x 0 0 32 0 INPUT NODEFVAL "data28x[31..0]"
-- Retrieval info: USED_PORT: data29x 0 0 32 0 INPUT NODEFVAL "data29x[31..0]"
-- Retrieval info: USED_PORT: data2x 0 0 32 0 INPUT NODEFVAL "data2x[31..0]"
-- Retrieval info: USED_PORT: data30x 0 0 32 0 INPUT NODEFVAL "data30x[31..0]"
-- Retrieval info: USED_PORT: data31x 0 0 32 0 INPUT NODEFVAL "data31x[31..0]"
-- Retrieval info: USED_PORT: data3x 0 0 32 0 INPUT NODEFVAL "data3x[31..0]"
-- Retrieval info: USED_PORT: data4x 0 0 32 0 INPUT NODEFVAL "data4x[31..0]"
-- Retrieval info: USED_PORT: data5x 0 0 32 0 INPUT NODEFVAL "data5x[31..0]"
-- Retrieval info: USED_PORT: data6x 0 0 32 0 INPUT NODEFVAL "data6x[31..0]"
-- Retrieval info: USED_PORT: data7x 0 0 32 0 INPUT NODEFVAL "data7x[31..0]"
-- Retrieval info: USED_PORT: data8x 0 0 32 0 INPUT NODEFVAL "data8x[31..0]"
-- Retrieval info: USED_PORT: data9x 0 0 32 0 INPUT NODEFVAL "data9x[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: USED_PORT: sel 0 0 5 0 INPUT NODEFVAL "sel[4..0]"
-- Retrieval info: CONNECT: @data 1 0 32 0 data0x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 10 32 0 data10x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 11 32 0 data11x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 12 32 0 data12x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 13 32 0 data13x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 14 32 0 data14x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 15 32 0 data15x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 16 32 0 data16x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 17 32 0 data17x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 18 32 0 data18x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 19 32 0 data19x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 1 32 0 data1x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 20 32 0 data20x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 21 32 0 data21x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 22 32 0 data22x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 23 32 0 data23x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 24 32 0 data24x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 25 32 0 data25x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 26 32 0 data26x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 27 32 0 data27x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 28 32 0 data28x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 29 32 0 data29x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 2 32 0 data2x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 30 32 0 data30x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 31 32 0 data31x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 3 32 0 data3x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 4 32 0 data4x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 5 32 0 data5x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 6 32 0 data6x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 7 32 0 data7x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 8 32 0 data8x 0 0 32 0
-- Retrieval info: CONNECT: @data 1 9 32 0 data9x 0 0 32 0
-- Retrieval info: CONNECT: @sel 0 0 5 0 sel 0 0 5 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux324.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux324.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux324.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux324.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL mux324_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
